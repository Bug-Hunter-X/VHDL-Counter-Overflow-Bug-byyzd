```vhdl
entity counter_fixed is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           count : out  integer range 0 to 7);
end entity;

architecture behavioral of counter_fixed is
    signal internal_count : integer range 0 to 7 := 0;
begin
    process (clk, rst)
    begin
        if rst = '1' then
            internal_count <= 0;
        elsif rising_edge(clk) then
            internal_count <= (internal_count + 1) mod 8; -- Modulo operation for wrap-around
        end if;
    end process;
    count <= internal_count; 
end architecture;
```